`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 06.02.2026 16:38:37
// Design Name: 
// Module Name: estimation_top
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module estimation_top (
    input  logic clk,
    input  logic reset,

    // tapped signals (read-only)
    input  logic pc_write,
    input  logic reg_write,
    input  logic mem_write,
    input  logic recovery_active
);


endmodule
